package my_package;

import uvm_pkg::*;

// UVM files
`include "uvm_macros.svh"
`include "my_sequence.sv"
`include "my_monitor.sv"
`include "my_driver.sv"
`include "my_agent.sv"
`include "my_scoreboard.sv"
`include "my_env.sv"
`include "my_test.sv"

endpackage
